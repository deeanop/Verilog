`timescale 1 ns/1 ps
module multiplexer4_to_1_tb;
	reg D0, D1, D2, D3, S0, S1;
	wire Y;
	multiplexer4_to_1 uut(
		.D0(D0),
		.D1(D1),
		.D2(D2),
		.D3(D3),
		.S0(S0),
		.S1(S1),
		.Y(Y)
	);
	initial begin
		$display("Time | D0 | D1 | D2 | D3 | S0 | S1 | Y");
		$monitor("%0t | %b | %b | %b | %b | %b | %b | %b ", $time, D0, D1, D2, D3, S0, S1, Y);
		S0 = 'b0; S1 = 'b0;
		D0 = 'b0; D1 = 'b0; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b1; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b1; D3 = 'b1; #10; 
		D0 = 'b1; D1 = 'b0; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b1; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b1; D3 = 'b1; #10;
		S0 = 'b0; S1 = 'b1;
		D0 = 'b0; D1 = 'b0; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b1; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b1; D3 = 'b1; #10; 
		D0 = 'b1; D1 = 'b0; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b1; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b1; D3 = 'b1; #10;
		S0 = 'b1; S1 = 'b0;
		D0 = 'b0; D1 = 'b0; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b1; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b1; D3 = 'b1; #10; 
		D0 = 'b1; D1 = 'b0; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b1; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b1; D3 = 'b1; #10;
		S0 = 'b1; S1 = 'b1;
		D0 = 'b0; D1 = 'b0; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b0; D2 = 'b1; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b0; D1 = 'b1; D2 = 'b1; D3 = 'b1; #10; 
		D0 = 'b1; D1 = 'b0; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b0; D2 = 'b1; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b0; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b0; D3 = 'b1; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b1; D3 = 'b0; #10;
		D0 = 'b1; D1 = 'b1; D2 = 'b1; D3 = 'b1; #10;
		$finish;
	end
endmodule		